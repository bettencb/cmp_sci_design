version https://git-lfs.github.com/spec/v1
oid sha256:0d47bbe25220e9336d36f5d71fd7adccb010d9e988306727e1457d9750d07097
size 4208
