version https://git-lfs.github.com/spec/v1
oid sha256:660dfca85fcc4c0dc8fc122891c57e42a260dc365e83378100ba3175d9b8e3ad
size 61583
