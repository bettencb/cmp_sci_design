version https://git-lfs.github.com/spec/v1
oid sha256:e26b9fb60d8a2ec8ab71506ef4807a308530e53862f7b146f46eca2a49af90e7
size 7824
