version https://git-lfs.github.com/spec/v1
oid sha256:a71cf6f8ceaa342772a4535ad02c1441c85779cc6814755dc8c419c4e55e14e0
size 11794
