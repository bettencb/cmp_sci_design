version https://git-lfs.github.com/spec/v1
oid sha256:ba8ffa1759a08c5fd304b28bf91ece521d34a147e9972e948acbf2bf55ba92fa
size 7920
