version https://git-lfs.github.com/spec/v1
oid sha256:7041d3a13ae8d12ab1f7e610e7293c8ab2f50c49f8dd57863dc70f187d9c7b48
size 12921
