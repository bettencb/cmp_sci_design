version https://git-lfs.github.com/spec/v1
oid sha256:7a5abdb681924a99c42631ab56b45e5f3817f5e797e903cba1d7ef5732c21a24
size 47660
