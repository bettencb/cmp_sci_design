version https://git-lfs.github.com/spec/v1
oid sha256:858fa0717ead39acbc4a6dc5735a67f833ec012bff3dfdd07c53894c536ed979
size 20997
