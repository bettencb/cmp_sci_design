version https://git-lfs.github.com/spec/v1
oid sha256:5f33d8fe15bc93676f0620b6138842355890618f05d1bee94173f51d2ef4e98a
size 48821
