version https://git-lfs.github.com/spec/v1
oid sha256:2f9e2c29edc4fbd39e282b04a3f05d0d35d591db5826b4a513b6026b01fc5e13
size 4075
