version https://git-lfs.github.com/spec/v1
oid sha256:9ada3d6ccea5e3f2cd15daa9cc0f22db9a3210a7a439df0d480e1d598b167e8b
size 5487
