version https://git-lfs.github.com/spec/v1
oid sha256:95de9b7617431ae3d825e018c0425a81efa6385a2ff5d46df8a236af9a500eca
size 16777
