version https://git-lfs.github.com/spec/v1
oid sha256:17e34b4f94a0edf657fd69d8e4c98d651e060da542015a7ded397720db2cb922
size 3792
