version https://git-lfs.github.com/spec/v1
oid sha256:fbb8b2b77f5bb652282e73ef23af5f759c938e80af7916f6e386805037286d48
size 11976
