version https://git-lfs.github.com/spec/v1
oid sha256:8cc67043432b6cedfa2ee6e2c2c5734aeaac8f4e4d7c5dcd991b0eca40fea1eb
size 8382
