version https://git-lfs.github.com/spec/v1
oid sha256:2bffa5b76fd27fce6af28a0d7d03dde79818567fcec5e68d3cbcd7fe6f89e096
size 7709
