version https://git-lfs.github.com/spec/v1
oid sha256:4986762116dc020201d713bf554225ae8a108c838f7f2faf30070ca94f0efbfa
size 8132
