version https://git-lfs.github.com/spec/v1
oid sha256:f05398a9b05e6fd6180b560e337cd377ded6c7fc1f6990147b1622d6f5c05328
size 8009
