version https://git-lfs.github.com/spec/v1
oid sha256:436c8c65b62e838febe5029a22b485c099f3ccd78c5810aaf71da682cbc2ddb8
size 66503
