version https://git-lfs.github.com/spec/v1
oid sha256:79d4ee432146c9ce3bf4863004214f930bccbfca80aebd5c08cbb4f857bac87b
size 4696
