version https://git-lfs.github.com/spec/v1
oid sha256:8b26d1954048605c5f6d830cc0c6c2e1eb93de4341851aff231f72c8cfb9f0ce
size 4844
