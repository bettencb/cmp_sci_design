version https://git-lfs.github.com/spec/v1
oid sha256:bffaa4a3c1459cca1413ad863b3a5e84d36e984af2c71b1a46416d330c5698f7
size 105726
