version https://git-lfs.github.com/spec/v1
oid sha256:fda8fa3792727403f5371c2ba67ab61fc1c0b0b1d14ddf39e812a591408fb3f4
size 2620
