version https://git-lfs.github.com/spec/v1
oid sha256:c52832d09a4cc4b0d2e748c22aca01553f2a05c3887d89387c9db5552f43535e
size 17249
