version https://git-lfs.github.com/spec/v1
oid sha256:f7348ee27d758bab7c3e34e09a847b26ee4242de14109f743070e2b674039897
size 3778
