version https://git-lfs.github.com/spec/v1
oid sha256:ac90ad5bd9406bacc335e87d6edeeb996983968b7eb5526e6306b14b7805ea95
size 3833
