version https://git-lfs.github.com/spec/v1
oid sha256:1c97a98ab8d7b05dc74cb1be755c4a80e288926d644d1b1b143b2a261f547f99
size 184859
