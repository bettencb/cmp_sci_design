version https://git-lfs.github.com/spec/v1
oid sha256:b2298eedda77bb1f52d1165ab7d609869d3b7c529acbe94ddeec316be9e1ee94
size 4684
