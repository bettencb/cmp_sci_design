version https://git-lfs.github.com/spec/v1
oid sha256:07d9467ece958cb64160dbf2897e071d65b930fda87975e223cd078efc0d7ed9
size 2620
