version https://git-lfs.github.com/spec/v1
oid sha256:0275635fda146340cd7ad74a41ff8b765381b7975f44a56663567c02dac668eb
size 3437
