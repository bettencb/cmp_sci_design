version https://git-lfs.github.com/spec/v1
oid sha256:f8efd65c3cc00d916a1a793ecac4d24c0418b2753f2c4b77adeb9c71cbcabc12
size 7940
