version https://git-lfs.github.com/spec/v1
oid sha256:1613977dabd6f75234ad5cd0afa3ba5cded96ceadc4e43eb064ae37a66eff91d
size 7719
