version https://git-lfs.github.com/spec/v1
oid sha256:c900b2311eaa4b09721649370378c9a1d46a667681ff5b88d98d05225119a2d9
size 5480
