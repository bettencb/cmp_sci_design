version https://git-lfs.github.com/spec/v1
oid sha256:a95676185f29946554a9db25a1334744e44b5545c93646e4d88c9c2ec285d128
size 3768
