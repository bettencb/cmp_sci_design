version https://git-lfs.github.com/spec/v1
oid sha256:3cc238bd36783cd51c132131addecb2ee7d6ffa9f29dc797f8e141b6a4ba5070
size 7564
