version https://git-lfs.github.com/spec/v1
oid sha256:e76e252730d5708bfef0e777cf634df7996452c75ca62e127c4830783540e244
size 25255
