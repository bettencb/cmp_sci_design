version https://git-lfs.github.com/spec/v1
oid sha256:9e82f563b52966f89f82c814be37150a917c9c98ac75020207e11461f785593a
size 14528
