version https://git-lfs.github.com/spec/v1
oid sha256:2df0c2b65cd6a351bada0d3bfb143e893b3599490bb0ecbb41c4b78e09eab02a
size 8216
