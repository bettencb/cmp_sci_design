version https://git-lfs.github.com/spec/v1
oid sha256:3e2e1cafe44b659a63e16810012e9fac257b153967302eac1f589ac315289b15
size 7316
