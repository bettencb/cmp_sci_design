version https://git-lfs.github.com/spec/v1
oid sha256:3bdfe2bba3b7d9857c85b34be298ab9c64a3d98835e27dfef518f321a806620b
size 13688
