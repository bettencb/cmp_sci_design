version https://git-lfs.github.com/spec/v1
oid sha256:1a6ea93ee6841857f2bb6201c955fa2071684b2cf7041e7a09863d1add312233
size 5485
