version https://git-lfs.github.com/spec/v1
oid sha256:764314fd8a7432898e88a47aae884a418f3c3d5bbd49e697022f7c972f67536a
size 3712
