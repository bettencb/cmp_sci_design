version https://git-lfs.github.com/spec/v1
oid sha256:fb34846cfdebc37cfeed748a751167df5df428554d73ea19a726849eb26eaae9
size 2733
