version https://git-lfs.github.com/spec/v1
oid sha256:578acd54ae86b1bc39bb643c45a6f0e276058182da6026e8f8e9044629c3077d
size 29991
