version https://git-lfs.github.com/spec/v1
oid sha256:44178b55a22c8d021f7a5632974a00cf3277e89a9908d40cfc349ab6c2b70215
size 7822
