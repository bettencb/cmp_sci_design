version https://git-lfs.github.com/spec/v1
oid sha256:e8b69cc38ca6c29bc0160f9a86357354382fc589642c9faedd27ea5953edf23b
size 4505
