version https://git-lfs.github.com/spec/v1
oid sha256:35dae8a7ee9619ee74c9baf6bc9c3b27d78a999ac03363161e4dd1ff9a1f6705
size 4676
