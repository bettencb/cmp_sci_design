version https://git-lfs.github.com/spec/v1
oid sha256:9bb4be235c269a0b7638652c65fee90ab2e7d46b7c18feb360f65f504e54d590
size 32226
