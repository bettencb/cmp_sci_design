version https://git-lfs.github.com/spec/v1
oid sha256:8a144f246bb6524fb85b48a69736b6de3fc89499d1d845372245f3ef629e1a0b
size 12923
