version https://git-lfs.github.com/spec/v1
oid sha256:2ec8d7ad3e40662bab3c968b0efd8cd96028eacebf417714acf735666ac62697
size 12132
