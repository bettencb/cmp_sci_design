version https://git-lfs.github.com/spec/v1
oid sha256:c25119f9c67d4655d9a9f934de5fbda5cf55a98f05d39b70e2d8b07f50fa09ef
size 4208
