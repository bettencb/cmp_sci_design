version https://git-lfs.github.com/spec/v1
oid sha256:7fff2d10638a77e11b1835f798ca05d8a50e8b52e8caf09db69c733c53356286
size 8463
