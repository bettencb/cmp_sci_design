version https://git-lfs.github.com/spec/v1
oid sha256:9d3feb68df8e2e6765f0f2041ba5917462feab842ce573560784faba776d0fef
size 5290
