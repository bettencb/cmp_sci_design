version https://git-lfs.github.com/spec/v1
oid sha256:210a9a3c8f133167b0070739f8c554848b583c95fa927854b420765d22e6ae3c
size 3459
