version https://git-lfs.github.com/spec/v1
oid sha256:95126ca0950a88c7487e4516a38f8402e7d1d03de9790fb76c0e913bf9ec8b32
size 7323
