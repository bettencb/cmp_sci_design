version https://git-lfs.github.com/spec/v1
oid sha256:df02a2139fc53e6bfec1529547422720a23f728078401cdae86429547ec3c4bb
size 4083
