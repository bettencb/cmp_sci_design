version https://git-lfs.github.com/spec/v1
oid sha256:0f213b5ac3037b939776717957b8463659723de2e977f3b9b1c755f6c51d4320
size 11113
