version https://git-lfs.github.com/spec/v1
oid sha256:6470ebc84aec7642f3dd787d6a8e39fd0da86adac49f4ce983160a9f64939714
size 30283
