version https://git-lfs.github.com/spec/v1
oid sha256:96006d96d8857941f870c58a6250bd3b42a480bc39c91f2ce5b0828c3c94ac26
size 8132
