version https://git-lfs.github.com/spec/v1
oid sha256:08aebf92648ba25ee5b4eb98643a76910d32d647b23fa95608860f502a0d34df
size 4855
