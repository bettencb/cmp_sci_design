version https://git-lfs.github.com/spec/v1
oid sha256:f200d98659708f08b7c86f3346c808229efd44e1d12f826771679b6c37196969
size 11328
