version https://git-lfs.github.com/spec/v1
oid sha256:2ad510298b5fea2167bf792d5c0e6bbfc62414fa24859a58c374027ba1c3ccb5
size 9351
