version https://git-lfs.github.com/spec/v1
oid sha256:9a1b32014b51239c085be0e1574577d06857603f970999461b656b2fa95b4ea3
size 8244
