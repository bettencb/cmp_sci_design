version https://git-lfs.github.com/spec/v1
oid sha256:c87855f419f1ec49f2307a5d06369b136e7c1a7df678b7c31b6625aeabd3b691
size 4693
