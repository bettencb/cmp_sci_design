version https://git-lfs.github.com/spec/v1
oid sha256:540bf7af7193d5392907a33cc829baf3eb41ebb17549923698e3d08478b097a8
size 8218
