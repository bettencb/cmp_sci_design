version https://git-lfs.github.com/spec/v1
oid sha256:8b19ae45c7ed2c0e5b4a4e278d99a3417366a9af369d28e1169804891eb0c807
size 3792
