version https://git-lfs.github.com/spec/v1
oid sha256:ac2fd60846a8748325c6291d39de9af38a7ba426b9b9dcf93feef36c44ab0c58
size 12126
