version https://git-lfs.github.com/spec/v1
oid sha256:b1afe4fdb03cb8c63ff985c7d48e4937fd8221b8dd8ef06f6a57281fe43b5152
size 7926
