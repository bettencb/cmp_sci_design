version https://git-lfs.github.com/spec/v1
oid sha256:b7c7f91ee924a547083b982e02a3e4acd059c364344c5a887e45cddf20c2014e
size 2892
