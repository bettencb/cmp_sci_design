version https://git-lfs.github.com/spec/v1
oid sha256:3139c43e42a9863fbb5e9e8e25945533fc5b40bb6d520b5f1f13ad695af4f830
size 8367
