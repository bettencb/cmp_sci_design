version https://git-lfs.github.com/spec/v1
oid sha256:02efd31f175789f2bb576a006df1c41295bd3f9b34136817c488e175ceb61c9e
size 7926
