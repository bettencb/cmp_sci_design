version https://git-lfs.github.com/spec/v1
oid sha256:b0c719ee30486e77cf6c354fdd9df142e5fcf3e7306f070ea1e889bda65f1273
size 8108
