version https://git-lfs.github.com/spec/v1
oid sha256:001bb41bc4ca630b7ed84725d877d19fabccb4242499383e1fe6aafd071aebdc
size 7866
