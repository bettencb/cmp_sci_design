version https://git-lfs.github.com/spec/v1
oid sha256:f3ebf3d46b551b43922e77650a58b997e147d8619f05018425dcdab361fa1750
size 3458
