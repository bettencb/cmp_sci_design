version https://git-lfs.github.com/spec/v1
oid sha256:d67662b7bb48b27dae7bae3c6fab7c602a010509393ab11ab0f4cdba042cc012
size 12535
