version https://git-lfs.github.com/spec/v1
oid sha256:731eae5a7edf7358dd80b75580772f35755d174d14c7db49721359984f616744
size 11387
