version https://git-lfs.github.com/spec/v1
oid sha256:dd7236815afb771740515653543a67d2280c4f0565e4d9605912546627791f8f
size 3019
