version https://git-lfs.github.com/spec/v1
oid sha256:f600c33d96705acefa5d8c853210b4f0249f9e52c3d269706974b4be41dbb5d2
size 8394
