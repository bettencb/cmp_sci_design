version https://git-lfs.github.com/spec/v1
oid sha256:d76c2918180a2221737034b82efcf5247dd636f433818133d856808ca4d1ff18
size 11043
