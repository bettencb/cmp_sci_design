version https://git-lfs.github.com/spec/v1
oid sha256:071803b5397d1b1d27afb25167a76e96ae291e06b66de9ce562e98071cf83671
size 2439
