version https://git-lfs.github.com/spec/v1
oid sha256:f7d7085e1282bb69df01148aca7cb70b595f4d12009de1c2f9eccb5d8179345e
size 22483
