version https://git-lfs.github.com/spec/v1
oid sha256:6a99f22cfb4b4ffe7b19cea1b55a439c1bc9cb33ef1406ff91cb1f96e156e5eb
size 6972
