version https://git-lfs.github.com/spec/v1
oid sha256:80b67f438e3a85900fcf65a2a0888a88643eee0fbb6570328e8f18ee5a3b4389
size 11761
