version https://git-lfs.github.com/spec/v1
oid sha256:8fe968b0eb14c6aef6ef7ad6ccfde6918752c410d7047115e5cf65aba8d4fc9b
size 10955
