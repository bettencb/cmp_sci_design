version https://git-lfs.github.com/spec/v1
oid sha256:5225f6c695f33d73226b65dda0b74bf7f7b704c90709f2571677ce18ea193f82
size 11578
