version https://git-lfs.github.com/spec/v1
oid sha256:4f0eb202612c81d2d0cfe83bd91d1c74f080d586711798deea5d5b531ada768d
size 11799
