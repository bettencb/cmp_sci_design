version https://git-lfs.github.com/spec/v1
oid sha256:41994affd2fbd593d45197939d3c55bb8c193eba1f545c862c49042e0840d807
size 16861
