version https://git-lfs.github.com/spec/v1
oid sha256:71d50ca03d0c65bab4ef0ee425fae1d2168ecede1ad1d2df5c2523f6607bbd31
size 7468
