version https://git-lfs.github.com/spec/v1
oid sha256:fa67aa83dc27de53a4cc3d907071c8eb97d3302efe78b05880a3fc89aeeaf7b8
size 8229
