version https://git-lfs.github.com/spec/v1
oid sha256:3dcc53c92a568396c991123233bcc317392dc0b3e1e97981885819fd071fe572
size 8306
