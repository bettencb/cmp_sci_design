version https://git-lfs.github.com/spec/v1
oid sha256:0b682a2eca506cfcca52d43f66c029490e0510c4bff6a2711530a4bb09e6c66b
size 7326
