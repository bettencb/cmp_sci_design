version https://git-lfs.github.com/spec/v1
oid sha256:e1db9b2d196a70ef5f822f246e33a9d1d837d4c93c954d591db20ff54081f532
size 7869
