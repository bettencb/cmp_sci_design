version https://git-lfs.github.com/spec/v1
oid sha256:32b24f0b50d6a02a44df00dac6894f1501342ec27171e6d236be43a2553805ea
size 3776
