version https://git-lfs.github.com/spec/v1
oid sha256:763222bfaad90fd060a2d4285804085e0712ea2ec5d44b82cc8b67f6318a3440
size 12065
