version https://git-lfs.github.com/spec/v1
oid sha256:27216a3dad93ab40d91e0d6b65b8066748acf1d1ace60c7d37230706244e2a38
size 12132
