version https://git-lfs.github.com/spec/v1
oid sha256:30940f8a62378fe0dbb9aaeda8a0e857646a0d2ada67ba706dd90fcffe395030
size 8052
