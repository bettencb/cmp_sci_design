version https://git-lfs.github.com/spec/v1
oid sha256:03fe2dbfb43eaf77f71978aaf7a37ff19d6dc48cb4d70f1a428b8d9ab00f47a4
size 22094
