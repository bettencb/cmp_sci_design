version https://git-lfs.github.com/spec/v1
oid sha256:d5cbe8a8cd3259481bfe673b2dd8b4f9063e9f47f52ea1c48b6cebe65f0d03b4
size 4697
