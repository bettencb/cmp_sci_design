version https://git-lfs.github.com/spec/v1
oid sha256:787b717f392f12a8c7479e80be6af7e50d7a6e453c5a30c8e5c7334fe8e0ee7f
size 11241
