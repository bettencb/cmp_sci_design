version https://git-lfs.github.com/spec/v1
oid sha256:c7611e20fec543ce79f4a88417ec70eaa72a284132e6049250b5b0bfe704446b
size 32226
