version https://git-lfs.github.com/spec/v1
oid sha256:e9a9838bcac7d43042ddf7f89d015859ecada591b533bb9f90d5b5c1bdb13691
size 5690
