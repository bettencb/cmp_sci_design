version https://git-lfs.github.com/spec/v1
oid sha256:b4726f3cf31c790926e1e761aadc6c76ebae1221bed62dd56ac1a2bffd5ff030
size 8497
