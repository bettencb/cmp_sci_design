version https://git-lfs.github.com/spec/v1
oid sha256:9601256865407c0f78db1bcf7ff1de5d0ee7843231a9612eed2469dd66470ec8
size 7473
