version https://git-lfs.github.com/spec/v1
oid sha256:717f7b9f6e34a7c40ad9ecbfc92e0499000513c213d464b323c2cad0aa6bdde4
size 3786
