version https://git-lfs.github.com/spec/v1
oid sha256:7d87f28a6e0cc6d1dc26cf711909ceea253615a53a36a89738a56b903920e820
size 7564
