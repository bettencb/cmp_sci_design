version https://git-lfs.github.com/spec/v1
oid sha256:4e4fcc1e33db2449bfbd93839495a2f382f82540cb1a4eb7d356e63f6511932b
size 1915296
