version https://git-lfs.github.com/spec/v1
oid sha256:95c5a54c144c4bdab000877bd4a180008e372aa5827a856d11550597da001222
size 3113
