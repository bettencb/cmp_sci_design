version https://git-lfs.github.com/spec/v1
oid sha256:9e90457622b8be8f8862cb47e801780413d5fca225a719ec4cba3f932e55efb6
size 11066
