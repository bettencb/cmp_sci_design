version https://git-lfs.github.com/spec/v1
oid sha256:ec6a6966164821d4b1b22edeec2eb5bd74fafede7bb582e0fdb495411cc3b6de
size 7648
