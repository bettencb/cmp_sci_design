version https://git-lfs.github.com/spec/v1
oid sha256:222929756c48c45e6c902da68472cf9462b334b42acf37fbcefec5b0fb13d4da
size 4685
