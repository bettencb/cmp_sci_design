version https://git-lfs.github.com/spec/v1
oid sha256:2babd117f7b4f0f4b7cf850e1f177e45685c3e0c9cbfdbd3e8ddfaaf989a43f2
size 8105
