version https://git-lfs.github.com/spec/v1
oid sha256:5f7621b73c6a94b04bc5f6aff98f91d56b7bc252e6ebb857107921fcb7ff9586
size 11387
