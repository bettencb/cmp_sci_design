version https://git-lfs.github.com/spec/v1
oid sha256:3d663a84ceed362aba3ba93eeaf387a9b705268c43322801dec7643e87ff91ff
size 7648
