version https://git-lfs.github.com/spec/v1
oid sha256:c5fdff178286b0778a5920e8a80a4bc5cccce276fdb2964072fbf1b34b94ff79
size 4216
