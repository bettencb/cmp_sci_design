version https://git-lfs.github.com/spec/v1
oid sha256:116969b584ee4f74b2f8dff53b0771b79b80eba921eff34efe3239e94a5dbe3e
size 7648
