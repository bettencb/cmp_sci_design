version https://git-lfs.github.com/spec/v1
oid sha256:c4b24b11377928ddd72415d01cf878a38f3674d77f9679fc94bc8cd404255177
size 4844
