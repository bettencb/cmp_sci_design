version https://git-lfs.github.com/spec/v1
oid sha256:254364d3f4de6a063ae87e5a04216b2bd6b1977e07f164bb9d4b05a8f68c4985
size 12123
