version https://git-lfs.github.com/spec/v1
oid sha256:6c921a9ef2874c5cbbcca63a14d2db95a363556a3497347ac0d1b359ab010c12
size 3704
