version https://git-lfs.github.com/spec/v1
oid sha256:9e22982c88fee3aeaf6cb49968896c46c2bcd8c4be09e6701fbc9bceefb34e5a
size 1676
