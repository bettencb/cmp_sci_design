version https://git-lfs.github.com/spec/v1
oid sha256:aa3bb84d71b5bb94fcb5795213216341bb0bbe8b273bc7b62905d41d2d938179
size 100722
