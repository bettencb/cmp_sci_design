version https://git-lfs.github.com/spec/v1
oid sha256:f341d9d2912509051d94090c63b093fbc7ac3c04de41c7a0dabb23627789aacd
size 11381
