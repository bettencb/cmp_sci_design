version https://git-lfs.github.com/spec/v1
oid sha256:3d11aec36aecf65a72f49edb0de302467eb7e1acc7c05d3e49b4207329411050
size 8660
