version https://git-lfs.github.com/spec/v1
oid sha256:21473709e3fb9db2b1552405e5fe82dced3fd1f329aad880ce762e588a35ddaa
size 3706
