version https://git-lfs.github.com/spec/v1
oid sha256:fd0195363456f22a8a0b49592184b00154b458a71278b81bbda81ce2798c5263
size 3818
