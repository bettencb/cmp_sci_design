version https://git-lfs.github.com/spec/v1
oid sha256:4c433d5051a4747a5ccac06d523ad96324b0cee30d52945c54e6ec22d16d24e3
size 3789
