version https://git-lfs.github.com/spec/v1
oid sha256:40e12faf1fcb6c7d5a353f131d66b3bb1d2b980e7d4673789a779db76bf43405
size 23294
