version https://git-lfs.github.com/spec/v1
oid sha256:36ae7382a7a1f64796ff05d68ac7c6a79d33daa5c27e510c528226e63cc9e30c
size 3019
