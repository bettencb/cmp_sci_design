version https://git-lfs.github.com/spec/v1
oid sha256:65a00861014875e9d1fdd6d00581fec0b2cdf6d8f7ce62cf5c1a81cd8cbe0aca
size 7734
