version https://git-lfs.github.com/spec/v1
oid sha256:6927ce8a8b9f561c9179e68a31bf6045eb9815090b86defaf9f25b10737d263c
size 4216
