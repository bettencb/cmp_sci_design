version https://git-lfs.github.com/spec/v1
oid sha256:7c877a8c8fa06e1b9dff40fdebd14e84f9705ed3b87fa04e4fb1776c3360c9f7
size 11787
