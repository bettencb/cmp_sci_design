version https://git-lfs.github.com/spec/v1
oid sha256:158928881ec7911323bfa6f855abc50ba06d5ecc22314774adef55d5cc9ff788
size 8327
