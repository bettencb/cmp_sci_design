version https://git-lfs.github.com/spec/v1
oid sha256:597033fde6a6600a5e51bafc2f7369aa39f01741c826f6c4510f3629f33d3afc
size 57032
