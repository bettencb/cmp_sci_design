version https://git-lfs.github.com/spec/v1
oid sha256:075309a4e30577a286c392503e51c6ec01aaf889bf61c55fdd0a9759b4f51777
size 10559
