version https://git-lfs.github.com/spec/v1
oid sha256:cc0f2561d297e3e76bcdc87bffd94bf8b2adf9dfe52f61642bfe41b3802e9220
size 4069
