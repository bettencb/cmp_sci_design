version https://git-lfs.github.com/spec/v1
oid sha256:9b69cba2f09b6c0c735246b9bca81bc3944869b330e8cf09fb69eabb2cfc0f91
size 1766
