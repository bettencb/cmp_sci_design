version https://git-lfs.github.com/spec/v1
oid sha256:fe589892288c8c4ba8d2133ebf32ee2a73c791fc5cea3a57ef191adafec348ac
size 8431
