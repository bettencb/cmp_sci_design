version https://git-lfs.github.com/spec/v1
oid sha256:d17f4770b85d3039af16f05ce15141a37c57b38c1511fef3b0cd32c8483ed6b1
size 4049
