version https://git-lfs.github.com/spec/v1
oid sha256:124d5dde3192f593bbdfb414d799f03b478b57d496e212988c5f1b97a1c72e69
size 5336
