version https://git-lfs.github.com/spec/v1
oid sha256:4fc05fb9a87743e6229501edfc288300435baa1660015262ee6efd913a20dbbe
size 7833
