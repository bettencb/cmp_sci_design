version https://git-lfs.github.com/spec/v1
oid sha256:9f66c7a794eef2b0145a0cd5d87588f9b220cea6148879907a94193dfb271a74
size 3464
