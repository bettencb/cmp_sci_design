version https://git-lfs.github.com/spec/v1
oid sha256:2b091fa8515c183fe9a89b6c0c2602fbc83649b02a5d6667cd403e8b5e001695
size 8132
