version https://git-lfs.github.com/spec/v1
oid sha256:aa0743523429bd3f3f355c454ae657aee298bd6fd3af1ca504e31db0b0128fd9
size 94004
