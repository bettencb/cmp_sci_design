version https://git-lfs.github.com/spec/v1
oid sha256:2da7818c7c84d20be7072d79788ba8b261e46073d98766806fc3ba9d9e980e2e
size 8756
