version https://git-lfs.github.com/spec/v1
oid sha256:335e1d89493b90a465b8394c068272f7c1b16ad73a4a9d38a336840be7dd7d77
size 11794
