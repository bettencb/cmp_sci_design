version https://git-lfs.github.com/spec/v1
oid sha256:0eef753e7ae71877f1cd63d8ce9c7defe34aa504254e894e5e1ddfb54042dd1f
size 3049
