version https://git-lfs.github.com/spec/v1
oid sha256:20964206f37c38c99f02ddb87a9a9f501703b3462c21455db989bc08907e221e
size 58227
