version https://git-lfs.github.com/spec/v1
oid sha256:88415f13e507f6511f7a72f6e41a40b82f5947a652d5604f797ae10f7a1fa808
size 11051
