version https://git-lfs.github.com/spec/v1
oid sha256:debde3736a090fb13824960b9189e6df603d1fe72fc6819ec10c69aea9a4a6e8
size 13711
