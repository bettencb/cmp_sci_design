version https://git-lfs.github.com/spec/v1
oid sha256:f76a75b47010d811f55758bce209868c191a3bee8807d87edc96be16f69591b3
size 4071
