version https://git-lfs.github.com/spec/v1
oid sha256:3d8380bf8a99e2ec808459605f84d17b1efe65386dce08347379ba3d9afa8893
size 20448
