version https://git-lfs.github.com/spec/v1
oid sha256:22044969938e470571b2d6f7178886ed250ff96999e644a5dbed51bbe0fd9d9a
size 12157
