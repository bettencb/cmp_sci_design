version https://git-lfs.github.com/spec/v1
oid sha256:6f86a666eeeb4f92342ee617c7223eafa068f97664972b1507eeba0d4fe62f09
size 43579
