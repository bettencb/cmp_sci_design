version https://git-lfs.github.com/spec/v1
oid sha256:9d3ecab6ab6e5818bc9b273d67cd9ce3d67dce2823aa2154e815f173df127532
size 9743
