version https://git-lfs.github.com/spec/v1
oid sha256:7ca2f414fffd21a4e9d610ec89955050eaf0cc5e1b41215ac9da82f466559a2c
size 6116
