version https://git-lfs.github.com/spec/v1
oid sha256:70ad014dbc83b574b92c79c596a4c2faa1eca68355c6a9aadb2cedd190af3522
size 23179
