version https://git-lfs.github.com/spec/v1
oid sha256:6eb3bb708d2ba642713f4179fa470ec553c6cf436f90bfd484ebe31e24e61b4b
size 8306
