version https://git-lfs.github.com/spec/v1
oid sha256:04fd98ac56c4f298904e84005672de40bb48c3181fc9ba69cadb88697f414b2d
size 66501
