version https://git-lfs.github.com/spec/v1
oid sha256:db0767b7c307d891efa1fd63b3c9e47667f1725c30868921fc47dc4a05ce0af2
size 5315
