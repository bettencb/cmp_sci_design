version https://git-lfs.github.com/spec/v1
oid sha256:a7c2f1c9c8fca7af2ae6373ca3960663ba0a484aac39114f763adbfc629b7c9c
size 3786
