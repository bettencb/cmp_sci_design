version https://git-lfs.github.com/spec/v1
oid sha256:b4f638d27a3f0948acd0d883183c5707202aff37a3017639f4908383e0206bb8
size 10376
