version https://git-lfs.github.com/spec/v1
oid sha256:a8d13a3be70a9fef3fa1f6cf60f2779a11609d947632ac313a8e3d573256d693
size 3438
