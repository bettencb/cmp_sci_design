version https://git-lfs.github.com/spec/v1
oid sha256:5ad5ae1081f05627eb51a46c305f0d596cbd1731511403c418136c3f639f83b1
size 4077
