version https://git-lfs.github.com/spec/v1
oid sha256:32fe76216254f478849969031277476b52001dca24c8e9d758d5aa52197e3de4
size 8209
