version https://git-lfs.github.com/spec/v1
oid sha256:ce7a01effaa8c9eb375fcdf97470761666e038e3e9a713b7c04f39326a1439d4
size 3828
