version https://git-lfs.github.com/spec/v1
oid sha256:91251b7088c81ff1856796e9bfa41a0d4b55bc2cca94911dae607f4cb96eb418
size 14467
