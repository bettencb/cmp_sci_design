version https://git-lfs.github.com/spec/v1
oid sha256:214bce6b1efa9ed4ba25ee2d6cca7c9263ad18a8d692db093ef0a060d25dfd44
size 20447
