version https://git-lfs.github.com/spec/v1
oid sha256:9d43e1025a812091710c93b01b1e2af5ef03fde5e56895b82730025fbbd7a805
size 29380
