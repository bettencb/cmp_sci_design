version https://git-lfs.github.com/spec/v1
oid sha256:ac18fffbeb9a55db40a5762078f019ac2ca7425498cf8ea915b24ba37e086390
size 8660
