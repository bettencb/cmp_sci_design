version https://git-lfs.github.com/spec/v1
oid sha256:75547211a652c6d16e3a0f76428246ce4677fd788dd4be83173dea7e7c5e2406
size 11121
