version https://git-lfs.github.com/spec/v1
oid sha256:17f373812d73cdd4f15fce4f3047ef470daef523b286e4318cd4afe32feab8f3
size 3833
