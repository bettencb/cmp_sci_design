version https://git-lfs.github.com/spec/v1
oid sha256:6b50415b4f64b2952a738961fc916b5caf36425bbe9995718dc9574e1a1f670c
size 4855
