version https://git-lfs.github.com/spec/v1
oid sha256:6336a0e5da93c4af4313f3fe981941e067e3b7e7b30a70d73db918df3b041b09
size 22639
