version https://git-lfs.github.com/spec/v1
oid sha256:7a995d8edb7c32d9190481a491e619dc17a806582e8df2ebddc14b5097926d78
size 107605
