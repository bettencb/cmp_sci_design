version https://git-lfs.github.com/spec/v1
oid sha256:1ccd3e6f0957cf290ade837ba29ea499c2023e0f9ddc59cee3841b0a2d108632
size 12382
