version https://git-lfs.github.com/spec/v1
oid sha256:adec3b0b2a04050cca944b341b33026e1b30cc80c047af576b151a43f3cec989
size 8621
