version https://git-lfs.github.com/spec/v1
oid sha256:0546354992f2c0bb229f6fdab54236f181c8e82751577025ede2eae105ecd7d4
size 7709
