version https://git-lfs.github.com/spec/v1
oid sha256:18fffbd996d2f89d962d5b03bdaeaa56dd985393f0f5c972348190e29fa569e2
size 3443
