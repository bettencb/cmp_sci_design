version https://git-lfs.github.com/spec/v1
oid sha256:b3731a1038b403f092bdbe257a65bc059801bd96160318b8ed176384ccaf2efb
size 11183
