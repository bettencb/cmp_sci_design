version https://git-lfs.github.com/spec/v1
oid sha256:632493b02e066298fe0ba2dbef86362c81292ba366b598f3b6993070399c3a19
size 36316
