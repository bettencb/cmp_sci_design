version https://git-lfs.github.com/spec/v1
oid sha256:d5721e06b72b0a80143e12ab0c7ab43171e0fc7401efc7c514f688dde5e06288
size 2800
