version https://git-lfs.github.com/spec/v1
oid sha256:ce76463fe720eeecc26c78e1724561583bc04d5e85d3ee804e6be3a8461fc142
size 7724
