version https://git-lfs.github.com/spec/v1
oid sha256:8a99777eb8def51abd2cf44186a19ff31fc61d81a9364805fcbef1c91efea402
size 3352
