version https://git-lfs.github.com/spec/v1
oid sha256:b9b5496302d2150402b8660139ca4b726becd2c551c95018d649ef9a374ddc18
size 11180
