version https://git-lfs.github.com/spec/v1
oid sha256:e053d48f706e99f542897cd2edda9aa0cefcd997a61095296708de8d055d4b95
size 4078
