version https://git-lfs.github.com/spec/v1
oid sha256:fab73041325dc2c49de9c9a60e5fbb37ffb84537636e2bf45ceb9dbb1896ddab
size 4524
