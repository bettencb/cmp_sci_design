version https://git-lfs.github.com/spec/v1
oid sha256:5981bfa0b79caf7a0ba4961e49415bfd355622281d3fffc483a6dbe53bc5aae5
size 4844
