version https://git-lfs.github.com/spec/v1
oid sha256:685e64647f40914acc37871cd4ea67dadc62382b4a4428b0bb32786b4400c815
size 1626
