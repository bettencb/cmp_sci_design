version https://git-lfs.github.com/spec/v1
oid sha256:817f9108e9f339104ac368dcf492ecebee75de3d6817d0699560b8418c2393eb
size 8114
