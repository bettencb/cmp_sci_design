version https://git-lfs.github.com/spec/v1
oid sha256:9180c50a71edda866b0a912cc4ecf6ea1f184117a833e3b3dce04189d527084a
size 3797
