version https://git-lfs.github.com/spec/v1
oid sha256:66ecfc68d98118f1683d1ab2593b08aed7675a664e3f5d3f417927e740219a90
size 11765
