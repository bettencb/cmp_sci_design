version https://git-lfs.github.com/spec/v1
oid sha256:c5efdf21f4cc6418fa08b2b524e292a63b9b7d4f2ab58be09c2cc686722fc6ea
size 17047
