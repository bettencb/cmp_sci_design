version https://git-lfs.github.com/spec/v1
oid sha256:7913db46ca2956172545bd9bfcd316ceba83b19645af04f19a55eb079c5bb062
size 8414
