version https://git-lfs.github.com/spec/v1
oid sha256:ccfa033a4a9764ae8c503597d97ad4da2ea6101170b1b90d5b585ef9dcdb2215
size 4206
