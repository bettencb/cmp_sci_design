version https://git-lfs.github.com/spec/v1
oid sha256:c2b996d37ddd74848b39b790c41ab5407ea4a3519c38a611f5f0076fad74f74e
size 4505
