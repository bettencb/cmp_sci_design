version https://git-lfs.github.com/spec/v1
oid sha256:150c8c8fc3dbca0627b781cb2a1fb878329c6a2831f11aabe8c6b1bde9b652ab
size 12695
