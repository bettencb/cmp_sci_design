version https://git-lfs.github.com/spec/v1
oid sha256:17c94750d757eff6cf061c60c5426ea75a18e571ee75de3dc19719d46d0e2faa
size 10232
