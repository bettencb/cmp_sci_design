version https://git-lfs.github.com/spec/v1
oid sha256:5ad5dc389ce83d3eba63fc948f0ad3642c50f58f13dcd48c5b97dfb5ea6c2ea7
size 3833
