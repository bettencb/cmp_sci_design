version https://git-lfs.github.com/spec/v1
oid sha256:5ea8b44ef467c8af37a2f2ef1935f0f707890b5ed70cb301ce4893764ec69b3c
size 96424
