version https://git-lfs.github.com/spec/v1
oid sha256:f538a1d1e4206d2b8fdf02a66c46cec29254afc520805395a1b9b154da2c6a7d
size 37092
