version https://git-lfs.github.com/spec/v1
oid sha256:1d483a743e830dd169d582850728a14036f639adab0d94aadbfd4aeefff3fc50
size 4653
