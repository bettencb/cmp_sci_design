version https://git-lfs.github.com/spec/v1
oid sha256:6ca17a41d363fed768360a2bef1b7def720451a0be61c9e5a37cb9651bcd3abc
size 11802
