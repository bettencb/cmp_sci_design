version https://git-lfs.github.com/spec/v1
oid sha256:8f9b0885ce05bdabbc8f37a14bf12d5ffc2775d1026fc4a3c930ded0a55c07d1
size 8396
