version https://git-lfs.github.com/spec/v1
oid sha256:767a99f74a16eb61fffeb4819e0de37450ca2e3791a42dcc2dc823d68b1a6554
size 12313
