version https://git-lfs.github.com/spec/v1
oid sha256:603190a27f6349998614d0fe68bdde9ff5414383cfb68a1b1f92f8e60bff1cb0
size 3792
