version https://git-lfs.github.com/spec/v1
oid sha256:43e1e64374c78f4aa19e68505c73e6e969fe5ed4729df35c29a30571126f4282
size 12927
