version https://git-lfs.github.com/spec/v1
oid sha256:43207ad125b7a4449fdaf23df34c33365372f7ba70710df96b10d6491bfdeca4
size 17120
