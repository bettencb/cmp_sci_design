version https://git-lfs.github.com/spec/v1
oid sha256:07749b2449982189e1471adff1403541e249aabaaa75433643533c37914f1b26
size 6996
