version https://git-lfs.github.com/spec/v1
oid sha256:cc2dd972d2a03969ae69e027308d0431cc407f8479a031bffffe88424bee6c39
size 5445
