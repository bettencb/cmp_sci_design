version https://git-lfs.github.com/spec/v1
oid sha256:7d301a66f6c7df31fb96babdebedbb3e94c8d188bb36512d76f1fc659669e3af
size 3451
