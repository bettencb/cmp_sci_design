version https://git-lfs.github.com/spec/v1
oid sha256:b1b6e89445296f1e3ba228b7488e4780c254b48dff5625c4d0f0af11445beaec
size 10858
