version https://git-lfs.github.com/spec/v1
oid sha256:9c8dbd119a1d164bf76d52a9510e18f7716528824bfdb916f2e63e5a823b8228
size 11753
