version https://git-lfs.github.com/spec/v1
oid sha256:63f88a7a590c28a7da3163795c0754a8ea856bebfa2d200295a61cdc76eb3b97
size 4697
