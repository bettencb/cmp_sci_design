version https://git-lfs.github.com/spec/v1
oid sha256:c36ce76e546040b93793e77de6f0184f50e67148762d29cb4d01933cae2dbd0d
size 3717
