version https://git-lfs.github.com/spec/v1
oid sha256:f143134843d9fb4ecc73f9b9b61308053e70e05a56eeb8fd651954dae9f7b721
size 4072
