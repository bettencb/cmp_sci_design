version https://git-lfs.github.com/spec/v1
oid sha256:86801b6767b4b86674d59adcb4ecfc46b51c301b1277f994bbc0eafd29c65062
size 7842
