version https://git-lfs.github.com/spec/v1
oid sha256:f35e9ada29a10aad1d64fd9b6fa9e572b45bb1500b545f0b56c8c321a51c108a
size 3446
