version https://git-lfs.github.com/spec/v1
oid sha256:3142dfc48287727307f9e75c9635562029f823bd9ed546f1793eb2023aeb8a64
size 8212
