version https://git-lfs.github.com/spec/v1
oid sha256:7452e5e9a8d11500fbfb01420715ad3dafe7cc6175ec79d1db3bc8878a622b15
size 13253
