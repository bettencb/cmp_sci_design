version https://git-lfs.github.com/spec/v1
oid sha256:9b0c45a7084912fc9f1c30bb1d174bf97a7b400d27bdf5d28a81014bf91cee52
size 13168
