version https://git-lfs.github.com/spec/v1
oid sha256:f31d043b541dbece7af17a8be0883a2d21d5793379b0304984a091a8958d0449
size 8752
