version https://git-lfs.github.com/spec/v1
oid sha256:29925b25814429ddf81f25480b16d6ac898298db98d4e808b4b264cf7ef2ca64
size 3438
