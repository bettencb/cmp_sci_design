version https://git-lfs.github.com/spec/v1
oid sha256:f3b5582f4037b99cce2d572030f88345fcbac611f28ddd67733c1bfaff5b2d47
size 2901
