version https://git-lfs.github.com/spec/v1
oid sha256:9f3dc49a999848634d875b3648195f2a2effa3f3c919e512da95075267af27c4
size 16363
