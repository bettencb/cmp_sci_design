version https://git-lfs.github.com/spec/v1
oid sha256:80549ff27032342061a18b4eb1d55e573f0067e6e75c7530f9d488a760b01e35
size 12918
