version https://git-lfs.github.com/spec/v1
oid sha256:d1d843bd82c7da2997824e63e22776e712d7f3a615b36cc54e6703a44d5f13e3
size 6116
