version https://git-lfs.github.com/spec/v1
oid sha256:2332b50c69c693bd2b24db622f1489067efb73054d8bdcc585e097b6edb5ce76
size 12132
