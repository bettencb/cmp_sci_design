version https://git-lfs.github.com/spec/v1
oid sha256:603217bdfc4b64a05c9037d82a7c9e74a70715856a4b7f3233f3b8801c188be2
size 4092
