version https://git-lfs.github.com/spec/v1
oid sha256:331fb7fcd7bd1ce78e6079d6a11d997f15be5e4713d5e93cd72d963d12a656bb
size 42719
