version https://git-lfs.github.com/spec/v1
oid sha256:339b6173dc9e99acec3d46380a7428459126d83f964609a72ba3d3f74456dd76
size 16470
