version https://git-lfs.github.com/spec/v1
oid sha256:a9a60937e17b50c02097224fb2f9c5328cca18f9d37e1877536fd4dd6a16e69c
size 12132
