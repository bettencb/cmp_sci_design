version https://git-lfs.github.com/spec/v1
oid sha256:f1addeaa6e7b8075b9557ea5adcb73acc3fb2123c495f950cd1c812eaf134bb7
size 13299
