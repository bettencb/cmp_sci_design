version https://git-lfs.github.com/spec/v1
oid sha256:627d5e16a1fd01ba4e4228e04cedaef078c6a5ea29acd735ea8d4974233eada9
size 11043
