version https://git-lfs.github.com/spec/v1
oid sha256:f72a299e6f4d528dadbcd00f606e3a72154341610c5492394480646d1b8e17d5
size 9665
