version https://git-lfs.github.com/spec/v1
oid sha256:cf7b144d1afdf9e2682276e64c5b02c0ad4dd1618b00a48d47d1efe942fc2099
size 7822
