version https://git-lfs.github.com/spec/v1
oid sha256:a2d196e99616aa6818f00305895b5ad1ba1b8781b4f2a17fd62ea2278e23c47b
size 7176
