version https://git-lfs.github.com/spec/v1
oid sha256:2b19192c0335f059ab21ebfab5fc3c123c65dc5a0470538d89a041f4125781cd
size 8754
