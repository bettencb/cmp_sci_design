version https://git-lfs.github.com/spec/v1
oid sha256:6b81859a7c4fd42f02aadb51f72df47a2e4af1c9e748ac806270348175906b91
size 17229
