version https://git-lfs.github.com/spec/v1
oid sha256:978556e9ae9cc335a0b13faac9e178562f2c5d44fc72dd1d38e93f6b295f6d54
size 7734
