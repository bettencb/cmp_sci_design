version https://git-lfs.github.com/spec/v1
oid sha256:f9dcc72d13d16912e86f26534f6457a4678cc9fb1f09d9922899822880094bd9
size 2895
