version https://git-lfs.github.com/spec/v1
oid sha256:ec391e4757ad63e9e4b1940af0cb46798eccbf20550bdf00762db0198f16ce28
size 7826
