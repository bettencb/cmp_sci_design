version https://git-lfs.github.com/spec/v1
oid sha256:016141ee4b8d7e9d8798fa0a9350e019945d05b6bf807206f98f1d2fede249ec
size 3309
