version https://git-lfs.github.com/spec/v1
oid sha256:95fd3a3550daad800b7018154d7609588fee7108dbfd7b05d06b72f6bca02e1a
size 4208
