version https://git-lfs.github.com/spec/v1
oid sha256:450f6e22647c99978ce27babaf5448b38e306057bedcb5585d1d4f5366ef358c
size 4069
