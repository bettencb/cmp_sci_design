version https://git-lfs.github.com/spec/v1
oid sha256:e42a319e7ea6ab8e39913cbac2d6e51884eff97168b9091b4c6653aa9b32a69a
size 7812
