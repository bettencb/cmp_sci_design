version https://git-lfs.github.com/spec/v1
oid sha256:5057af8700b380f4d61bf328e89a9c6e7648496830870c13021cf7a6644a3c53
size 12926
