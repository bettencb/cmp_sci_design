version https://git-lfs.github.com/spec/v1
oid sha256:5170412bd98c248025b76d7baaae70e656a8d72a98b83383269aa9fb28f79dd1
size 7951
