version https://git-lfs.github.com/spec/v1
oid sha256:f88a546009b2f6eb917aa84be81db7805468a8caa14a9f2df0b845ccf4178da3
size 4705
