version https://git-lfs.github.com/spec/v1
oid sha256:f1edd35f16997e3c66ae779275315379e1123d37878e25df4b6d670e1d845bc4
size 4201
