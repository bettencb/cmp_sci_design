version https://git-lfs.github.com/spec/v1
oid sha256:0c4bce62c824b41ba2b23f45a20fb58e160c3c4d5b02f85321ce26986a4935c0
size 7319
