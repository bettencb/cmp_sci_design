version https://git-lfs.github.com/spec/v1
oid sha256:361227ea9d27084185466ebdcb07d69fe043a034c11f629bbefa58d76cf59146
size 13291
