version https://git-lfs.github.com/spec/v1
oid sha256:188880d79a6cd5d25f100fbac6bb6fe3cea2a266dcf786c15edd7e0b9684caf9
size 61583
