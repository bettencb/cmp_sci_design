version https://git-lfs.github.com/spec/v1
oid sha256:2da5eb441efb864cd191bbb52ec01603dd12c39665ff3e989f6af4dd4ea4de9c
size 3572
