version https://git-lfs.github.com/spec/v1
oid sha256:538c21b2b3ffdbbfc96c9246f333c5ceffd9bab2c9ae535513730fe23ef6b45d
size 8309
