version https://git-lfs.github.com/spec/v1
oid sha256:3649f4343e47f0168ef8e931b15a3d4b3b371566d2659407384f6f631145a296
size 5610
