version https://git-lfs.github.com/spec/v1
oid sha256:20a199db2a31d54662fe25868422df21abcdb8eba626fa0e1fdd808036a8584e
size 7926
