version https://git-lfs.github.com/spec/v1
oid sha256:00100a70cdb92744426a2b203d3e30e401c77b38ef1efa83468dd790f4c992be
size 4208
