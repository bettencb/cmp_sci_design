version https://git-lfs.github.com/spec/v1
oid sha256:12a614f35dc04b68b93b0bfe4efd8ec3352086836701e2439de759555ca1777e
size 7648
