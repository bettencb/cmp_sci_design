version https://git-lfs.github.com/spec/v1
oid sha256:97627dd912881d2330d6eb39d40049af7db122b34e48129eaf6f5d9000b925c8
size 7564
