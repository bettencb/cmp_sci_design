version https://git-lfs.github.com/spec/v1
oid sha256:de3713087dde66d9780e53f1f722d2aeb735193d4b201f82854383b773afd2b8
size 5328
