version https://git-lfs.github.com/spec/v1
oid sha256:6f7b12710319f6a57df467c888219d5d18c036dcd1b52331fcb4386745eb3e89
size 3792
