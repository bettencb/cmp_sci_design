version https://git-lfs.github.com/spec/v1
oid sha256:b8dfd0b94fb2d5e859ed5da1b6d42e13c4cd7768d57cd500ce892855c746f820
size 3459
