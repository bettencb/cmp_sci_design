version https://git-lfs.github.com/spec/v1
oid sha256:af5f89c40aa88ef626395f2d739f4f3e13852e215dc6c82b591834e5a58497d0
size 7954
