version https://git-lfs.github.com/spec/v1
oid sha256:1e517b895f2a7684295aaf36f4a6c2b0e74a3d734ab5d6f5517e74887660f4c2
size 12157
