version https://git-lfs.github.com/spec/v1
oid sha256:b38fc5d1c46593f8146001ee0e46b90a318fb3d82935ccf47b7a78b9d36a99cb
size 8739
