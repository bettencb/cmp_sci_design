version https://git-lfs.github.com/spec/v1
oid sha256:98245e4a7875497ff67a6bf18c59a4d3128f9c8df82b893881c913445ba35046
size 7832
