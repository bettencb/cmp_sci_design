version https://git-lfs.github.com/spec/v1
oid sha256:8113f415b57f955e479c4467cec17514208fcc952aae02bccc1bfae823f5b26e
size 9519
