version https://git-lfs.github.com/spec/v1
oid sha256:01eb9771836d3331dee40f3e0c399512f57903a0b9d7499eeaf8130c70d3bc91
size 3797
