version https://git-lfs.github.com/spec/v1
oid sha256:b17e0a637f8839c0c40b7faeba4bfb2dfefbc4f8dddffb2795b3a59fd0b2d1d8
size 5379
