version https://git-lfs.github.com/spec/v1
oid sha256:5f51a9dc5594eeb629a0733212f7949bb68cf8d565326cd475d75cb9889c3f46
size 5962
