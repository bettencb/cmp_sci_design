version https://git-lfs.github.com/spec/v1
oid sha256:a0a95a09a9e319bb49544e6330267aaeff83d99429508d12e7555816f0690c70
size 119890
