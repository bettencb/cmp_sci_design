version https://git-lfs.github.com/spec/v1
oid sha256:2345f011bed4230c95ddf92290828ef4c92bf8886d13851a5c73c577bd0b3760
size 8122
