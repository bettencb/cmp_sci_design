version https://git-lfs.github.com/spec/v1
oid sha256:352df1fb2feb8ea73220fc191121422a87d2083e17cac5e7208f8b742e3c5946
size 8215
