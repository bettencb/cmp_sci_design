version https://git-lfs.github.com/spec/v1
oid sha256:9bdc1e8aaf6425e87461833efac1ffdb8d16de7d6eac6aaecf73465d5eded94c
size 33038
