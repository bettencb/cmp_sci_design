version https://git-lfs.github.com/spec/v1
oid sha256:e90604f2b68fb8ce931307a4b27ab3d203c1ac9b6280fabbba0efaae7a1c719f
size 9260
