version https://git-lfs.github.com/spec/v1
oid sha256:274bd655665f0c4ab335eedf2495a3570b4aada544ac9820fa7a17c1688a0bc9
size 8292
