version https://git-lfs.github.com/spec/v1
oid sha256:465e3b88c018ece9efcf735b008ce0b4ff6e15d4733cd38e0bf47884b8df0a07
size 7967
