version https://git-lfs.github.com/spec/v1
oid sha256:ee84544d343a599ab8305fe26f8a95996601fffceef9e73331ab59678c054f40
size 3465
