version https://git-lfs.github.com/spec/v1
oid sha256:8f371395198f28b49eefded5424946622187e1adb3c699ca2b60238d0c2c7813
size 182983
