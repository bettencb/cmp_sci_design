version https://git-lfs.github.com/spec/v1
oid sha256:062dc11412f82a311c1d1b9d5585903cb382dfe3bf8a9879b0f11b2420cf56ff
size 1633
