version https://git-lfs.github.com/spec/v1
oid sha256:06c877fa8704be270543f2edec7c8a94c5518f097981ec7a3b2ebe318801fb3a
size 119386
