version https://git-lfs.github.com/spec/v1
oid sha256:425d786cb1966a668fd48fbfee67af5eea7e83d8c7c5edeeeb8d9c7c633fb6d1
size 7974
