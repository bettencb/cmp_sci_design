version https://git-lfs.github.com/spec/v1
oid sha256:87bc169db89523e21869d5cc5a144b074731506da2a14cd3fa9e9a2f538a85fb
size 13697
