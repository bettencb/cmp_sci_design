version https://git-lfs.github.com/spec/v1
oid sha256:7a672547ea4016eb749a798fcc9372f9630a0a6098c158e4a94ac37ee4442e1d
size 3311
