version https://git-lfs.github.com/spec/v1
oid sha256:c0b9b06dd4d154e1d31d79273e27b2a0af1162100e2453d74620d5060d778816
size 12918
