version https://git-lfs.github.com/spec/v1
oid sha256:6cb2d8f13f7f7d337499d6d5d5468d45f3f3ed5f9658a4d63cdb2d9d5fc47cd3
size 42240
