version https://git-lfs.github.com/spec/v1
oid sha256:2c98949944714e4183a0bfe5ae1d96b3d2b2b624fabfe36901c10e99f5e3ea76
size 4103
