version https://git-lfs.github.com/spec/v1
oid sha256:e5233962c242013c2967be739a56289651f3c802c772a4a7249b14c23ab24abf
size 4208
