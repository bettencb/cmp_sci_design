version https://git-lfs.github.com/spec/v1
oid sha256:70dfb18ce7cd42bf7e8955fa7f643394a9ad1ff32bfc666a73f0bb06973cd7db
size 8493
