version https://git-lfs.github.com/spec/v1
oid sha256:3ea9483ede0bce9404f8abd0c8498fe9062198d45053ac7cdb48b960b245cbcd
size 7882
