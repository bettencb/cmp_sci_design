version https://git-lfs.github.com/spec/v1
oid sha256:1f84d054513e78e06f0de4dec7c8c39653ffcf1a3001f5467bedfbbe5f470987
size 8132
