version https://git-lfs.github.com/spec/v1
oid sha256:cc1136b226dff678bed2ec4b753005c45700140cc78b83267edab86590f150bc
size 17332
