version https://git-lfs.github.com/spec/v1
oid sha256:0061d5ee44d06a3e42bacc609086733633a6541d7500ad646170500e5cb2a12c
size 11387
