version https://git-lfs.github.com/spec/v1
oid sha256:c44de569e2bc513b9f8d9ec0401300857936d20beb56815e2536caea8b4c5492
size 11790
