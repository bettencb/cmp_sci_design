version https://git-lfs.github.com/spec/v1
oid sha256:2f9f663eecde0c0acb002e8f1dc9cd7364875d4759eed3d743cdd0c00449a14b
size 13697
