version https://git-lfs.github.com/spec/v1
oid sha256:4229e99d2d8cd8a9c9cac6ebdedf1e7c26a18671f170ea38cd9ae1b6ab1bc00a
size 31042
