version https://git-lfs.github.com/spec/v1
oid sha256:42d1f6d4370a89dec6f99889220155c020b118c8a9ce7a0b3bc0e34df071c39c
size 3737
