version https://git-lfs.github.com/spec/v1
oid sha256:f7299cc9c06bec3a97670c77f341b0f43b7d223a09b20e568391a0c01fbb227d
size 4501
