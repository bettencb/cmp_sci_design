version https://git-lfs.github.com/spec/v1
oid sha256:9a0a6133a79d5b4126106fc9cc62009e8ded8ac5f1a11e913e03ae1cf1d197a0
size 8195
