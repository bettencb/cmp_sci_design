version https://git-lfs.github.com/spec/v1
oid sha256:aad6fcd88ff9de2c294a5ce3db4c124f418938f3e2dd2f289b319f070c609216
size 7316
