version https://git-lfs.github.com/spec/v1
oid sha256:6a82716da4a2fc74ba422f0a7156fcfa9777951201effe2ed90ec16714281134
size 16006
