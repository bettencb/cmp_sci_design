version https://git-lfs.github.com/spec/v1
oid sha256:365b817ff5f491472387606b951a350d8242025a64fb4bb6b9480afe5ee1ce09
size 13426
