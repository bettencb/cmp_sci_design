version https://git-lfs.github.com/spec/v1
oid sha256:e6886972d7b016116cbb01f706dd0e7481a112ca7b78775beb13a969a43251a5
size 2641
