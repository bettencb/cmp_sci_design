version https://git-lfs.github.com/spec/v1
oid sha256:71884b63e9f8f1cbdd2cb7f0d01a061384dec4fdb3b432fbca093553ec69ac5c
size 7926
