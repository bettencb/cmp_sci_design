version https://git-lfs.github.com/spec/v1
oid sha256:8ed88c55d0080b872c82b3f4cc2a329431905bc9742e43e98fa8a14d2e6fd7b8
size 11773
