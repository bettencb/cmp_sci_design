version https://git-lfs.github.com/spec/v1
oid sha256:dfe5eb0473125e651ce707140be38c3284cf25c4e295ac5c554708b43c300c94
size 3572
