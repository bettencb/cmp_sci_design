version https://git-lfs.github.com/spec/v1
oid sha256:8b3395a496903c6af787defdd6a084462784a6ba2446e9e07124ece84886bd38
size 8493
