version https://git-lfs.github.com/spec/v1
oid sha256:0de4814973335211aa89ccee9e8699583403b007ceb6d86750a17d1c73c0e6ce
size 3637
