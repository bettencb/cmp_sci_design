version https://git-lfs.github.com/spec/v1
oid sha256:e5a14ce16f40262d653ba96d8bbd4f43363db0206d12fc1ee3075b92f735aca9
size 4028
