version https://git-lfs.github.com/spec/v1
oid sha256:fef02a95faa3ef52884222f3e00e466794799660a58ff7bb9e7a63ecfc8e8f89
size 11797
