version https://git-lfs.github.com/spec/v1
oid sha256:e501871079decc606a6c160977a8b78c4f23801ebbc6cea11633a5d32e72b593
size 3701
