version https://git-lfs.github.com/spec/v1
oid sha256:90846cb9af6a52de4fd87331c36fb69185c47d2357d3dd8de32a36b11b2223fa
size 12157
