version https://git-lfs.github.com/spec/v1
oid sha256:2943ef61abc52798bc17f21852e6ff2c1a7e046e608d6cb602b65f03e67b94f5
size 6103
