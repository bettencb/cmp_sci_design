version https://git-lfs.github.com/spec/v1
oid sha256:90ece6394c3ccb478f8bd70b3d98b27a468c4d5fba9d131db183a7e580f7fa6c
size 11358
