version https://git-lfs.github.com/spec/v1
oid sha256:c73eb40d96c36a159de0c395a5f2c077800bee90f0d2700cd84802aa275c4692
size 8396
