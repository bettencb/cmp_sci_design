version https://git-lfs.github.com/spec/v1
oid sha256:1ef14931a15742bf1722ee08d3acf17c7b0d06375c62ff4d1539e197d35d8a17
size 6752
