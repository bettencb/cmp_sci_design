version https://git-lfs.github.com/spec/v1
oid sha256:46cae06b6ec44e9c57757d3889cdc2b1089c063b820a1e84853d027a404f1888
size 3664
