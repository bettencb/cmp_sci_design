version https://git-lfs.github.com/spec/v1
oid sha256:240e5df7bf217b6ec354e0585b3f61677f2d3896629fb22ec1c6babd2dd72ec0
size 7458
