version https://git-lfs.github.com/spec/v1
oid sha256:802464660dfbd22cdfb3a2eac0dc63b4ad0d534a55889269e83c8468aa63942c
size 3724
