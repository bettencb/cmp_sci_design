version https://git-lfs.github.com/spec/v1
oid sha256:03dc261285c91781ba5d90831266afc3aeda28878fd6e657acff4c7c61d6608d
size 7857
