version https://git-lfs.github.com/spec/v1
oid sha256:5187044e34f47fb42fc17a1820a290fd43542866cc9961ba5ee0b1aa77210127
size 16777
