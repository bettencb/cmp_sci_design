version https://git-lfs.github.com/spec/v1
oid sha256:97e7d91ef3654ba3c1dac747da1026141734120faeeee761f1fd40c7b5f2ccc6
size 4524
