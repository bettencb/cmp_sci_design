version https://git-lfs.github.com/spec/v1
oid sha256:5caa79e6e38ced76045ae2dd04109bf13392fb893c28691f05869139235a42ea
size 6146
