version https://git-lfs.github.com/spec/v1
oid sha256:8d62f728c03f2c590ac1ed3eb622917f31372bd0be2032b8ca85e47735cc55d6
size 7150
