version https://git-lfs.github.com/spec/v1
oid sha256:498028efe22216dd1c233a8d31c736a9fc276b9148ab27808d842d9fc553e5db
size 16334
