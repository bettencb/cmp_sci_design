version https://git-lfs.github.com/spec/v1
oid sha256:18441e95d19657e2d637c64f4756af80997aae0b408d48cfea087cee3168762f
size 4855
