version https://git-lfs.github.com/spec/v1
oid sha256:660edfa8e8c559f378108a271252f68ae416bf53b0478714f1d49fe6b6005150
size 3828
