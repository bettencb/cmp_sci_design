version https://git-lfs.github.com/spec/v1
oid sha256:58d7be8ad29e1d8526e995651ba9d07ac8e6f5f2bd699641bde0a3a5296d6309
size 3350
