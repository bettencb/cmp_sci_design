version https://git-lfs.github.com/spec/v1
oid sha256:bb1f5a98f351853246cad0105422098816e5eb1e7d3551272e1c42cd5b075e82
size 11045
